
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY OrGate IS
    PORT(
        i_a : IN STD_LOGIC_VECTOR(3 downto 0);
i_b : IN STD_LOGIC_VECTOR(3 downto 0);

        o_a : OUT STD_LOGIC_VECTOR(4 downto 0);

    );
END OrGate;

ARCHITECTURE behavioral_OrGate OF OrGate IS
BEGIN

END behavioral_OrGate;
